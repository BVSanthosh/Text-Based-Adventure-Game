bedroom
[("bedroom",Room {room_desc = "You are in your bedroom.", exits = [Exit {exit_dir = North, exit_desc = "To the north is a kitchen. ", room = "kitchen"}], objects = [Obj {obj_name = "mug", obj_longname = "a coffee mug", obj_desc = "A coffee mug", isHeavy = False}]}),("kitchen",Room {room_desc = "You are in the kitchen. The back door is closed.", exits = [Exit {exit_dir = South, exit_desc = "To the south is your bedroom. ", room = "bedroom"},Exit {exit_dir = East, exit_desc = "To the east is a hallway. ", room = "hall"}], objects = [Obj {obj_name = "cupboard", obj_longname = "the cupboard you keep your coffee pot in", obj_desc = "The cupboard is locked.", isHeavy = True}]}),("hall",Room {room_desc = "You are in the hallway. The front door is closed. The basement door is locked.", exits = [Exit {exit_dir = North, exit_desc = "To the north is the front door. ", room = "locked"},Exit {exit_dir = West, exit_desc = "To the west is a kitchen. ", room = "kitchen"},Exit {exit_dir = East, exit_desc = "To the east is the hallway extension. ", room = "hall extension"},Exit {exit_dir = South, exit_desc = "To the south is the door to the basement. ", room = "locked"}], objects = []}),("street",Room {room_desc = "You have made it out of the house.", exits = [Exit {exit_dir = In, exit_desc = "You can go back inside if you like. ", room = "hall"}], objects = []}),("hall extension",Room {room_desc = "You are in the later part of the hallway.", exits = [Exit {exit_dir = West, exit_desc = "To the west is the main hallway. ", room = "hall"},Exit {exit_dir = North, exit_desc = "To the north is a useless room. ", room = "useless"},Exit {exit_dir = East, exit_desc = "To the east is a useless room. ", room = "useless"},Exit {exit_dir = South, exit_desc = "To the south is the diner. ", room = "diner"}], objects = []}),("diner",Room {room_desc = "You are in the diner.", exits = [Exit {exit_dir = North, exit_desc = "To the north is the hallway.", room = "hall extension"}], objects = [Obj {obj_name = "tv", obj_longname = "a TV playing a video-tape", obj_desc = "The video-tape reminds you of the safe password!", isHeavy = True},Obj {obj_name = "safe", obj_longname = "a combination safe you keep your basement key in", obj_desc = "The safe is locked. You remember recording the password.", isHeavy = True},Obj {obj_name = "statue", obj_longname = "a broken statue holding something", obj_desc = "The kitchen cupboard key is stuck in the hands of the broken statue. If you fixed it you could get the key.", isHeavy = True}]}),("basement",Room {room_desc = "You are in the basement.", exits = [Exit {exit_dir = North, exit_desc = "To the north is the stairs to hallway.", room = "hall"}], objects = [Obj {obj_name = "hand", obj_longname = "a stone hand", obj_desc = "A stone hand that looks similar to the other one on the statue in your diner.", isHeavy = False},Obj {obj_name = "beans", obj_longname = "fresh coffee beans", obj_desc = "The coffee beans you store in the basement. Luckily you already brewed a pot this morning and left it in the cupboard.", isHeavy = False},Obj {obj_name = "monster", obj_longname = "a big, angry monster that glares when you get too close", obj_desc = "When you try get a closer look at it, the monster suddenly growls and lunges at you! You have died!", isHeavy = True}]})]
[]
False
False
False
False
False